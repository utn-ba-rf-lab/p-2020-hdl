
// ASCII Characters
	parameter U_ASCII = 8'd85;
	parameter T_ASCII = 8'd84;
	parameter N_ASCII = 8'd78;
	parameter O_ASCII = 8'd79;
	parameter K_ASCII = 8'd75;
	parameter E_ASCII = 8'd69;
	parameter R_ASCII = 8'd82;
	parameter v_ASCII = 8'd118;
	parameter _2_ASCII = 8'd50;

// Samp Rates
	parameter SAMP_RATE_8K 	 = 16'd8000;
	parameter SAMP_RATE_11K  = 16'd11025; // 11.025k
	parameter SAMP_RATE_16K  = 16'd16000;
	parameter SAMP_RATE_22K  = 16'd22050; // 22.05k
	parameter SAMP_RATE_24K  = 16'd24000;
	parameter SAMP_RATE_32K  = 16'd32000;
	parameter SAMP_RATE_44K  = 16'd44100; // 44.1k
	parameter SAMP_RATE_48K  = 16'd48000;
	parameter SAMP_RATE_0K   = 16'd0;

// FSM STATES
	parameter ST_0   = 5'd0;
	parameter ST_1   = 5'd1;
	parameter ST_2   = 5'd2;
	parameter ST_3   = 5'd3;
	parameter ST_4   = 5'd4;
	parameter ST_5   = 5'd5;
	parameter ST_6   = 5'd6;
	parameter ST_7   = 5'd7;
	parameter ST_8   = 5'd8;
	parameter ST_9   = 5'd9;
	parameter ST_10  = 5'd10;
	parameter ST_11  = 5'd11;
	parameter ST_12  = 5'd12;
	parameter ST_13  = 5'd13;
	parameter ST_14  = 5'd14;
	parameter ST_15  = 5'd15;
	parameter ST_16  = 5'd16;
	parameter ST_17  = 5'd17;
	parameter ST_18  = 5'd18;
	parameter ST_19  = 5'd19;
	parameter ST_20  = 5'd20;
